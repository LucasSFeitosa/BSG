module BSG(
	input logic [7:0]BSG_CONTROL,
	input logic [7:0]BSG_DATA_1,
	input logic [7:0]BSG_DATA_2,
	
	input SYS_CLK, G_CLK_TX, reset
);

//modulador modulador_h(.saida(), .dado(), .clk(G_CLK_TX), .reset(reset))


endmodule