//AMBA comunicaç~ao